`ifndef I2C_SCOREBOARD_SV
`define I2C_SCOREBOARD_SV

//==============================================================================
// I2C Scoreboard
//
// Professional scoreboard with:
// - TLM Analysis FIFO for decoupled processing
// - Expected vs Actual comparison
// - uvm_event integration for synchronization
// - uvm_callback hooks for extensibility
// - Statistical tracking and reporting
//==============================================================================

class i2c_scoreboard extends uvm_scoreboard;
  `uvm_component_utils(i2c_scoreboard)
  
  // Register callback type
  `uvm_register_cb(i2c_scoreboard, i2c_scoreboard_callback)
  
  //----------------------------------------------------------------------------
  // TLM Ports
  //----------------------------------------------------------------------------
  uvm_tlm_analysis_fifo #(i2c_transaction) analysis_fifo;
  uvm_analysis_imp #(i2c_transaction, i2c_scoreboard) item_imp;
  
  //----------------------------------------------------------------------------
  // Expected Transaction Queue
  //----------------------------------------------------------------------------
  i2c_transaction expected_queue[$];
  
  //----------------------------------------------------------------------------
  // Statistics
  //----------------------------------------------------------------------------
  int unsigned total_received  = 0;
  int unsigned total_compared  = 0;
  int unsigned total_matched   = 0;
  int unsigned total_mismatched = 0;
  
  //----------------------------------------------------------------------------
  // Configuration
  //----------------------------------------------------------------------------
  bit enable_comparison = 1;
  
  //----------------------------------------------------------------------------
  // Events for Synchronization
  //----------------------------------------------------------------------------
  uvm_event transaction_received_event;
  uvm_event comparison_done_event;
  uvm_event mismatch_event;
  
  //----------------------------------------------------------------------------
  // Constructor
  //----------------------------------------------------------------------------
  function new(string name, uvm_component parent);
    super.new(name, parent);
    item_imp = new("item_imp", this);
  endfunction
  
  //----------------------------------------------------------------------------
  // Build Phase
  //----------------------------------------------------------------------------
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    
    // Create TLM FIFO
    analysis_fifo = new("analysis_fifo", this);
    
    // Create events
    transaction_received_event = new("transaction_received_event");
    comparison_done_event = new("comparison_done_event");
    mismatch_event = new("mismatch_event");
    
    `uvm_info("SCB", "Scoreboard built with TLM FIFO and event synchronization", UVM_MEDIUM)
  endfunction
  
  //----------------------------------------------------------------------------
  // Write Function - Called by Monitor via Analysis Port
  //----------------------------------------------------------------------------
  function void write(i2c_transaction tr);
    i2c_transaction tr_copy;
    
    total_received++;
    
    // Clone transaction for FIFO
    tr_copy = i2c_transaction::type_id::create("tr_copy");
    tr_copy.copy(tr);
    
    // Push to FIFO for async processing
    analysis_fifo.write(tr_copy);
    
    // Trigger event
    transaction_received_event.trigger(tr_copy);
    
    `uvm_info("SCB", $sformatf("Received transaction #%0d: %s", 
              total_received, tr.convert2string()), UVM_HIGH)
  endfunction
  
  //----------------------------------------------------------------------------
  // Run Phase - Comparison Loop
  //----------------------------------------------------------------------------
  task run_phase(uvm_phase phase);
    i2c_transaction actual_tr;
    
    forever begin
      // Get transaction from FIFO (blocking)
      analysis_fifo.get(actual_tr);
      
      if (enable_comparison && expected_queue.size() > 0) begin
        compare_with_expected(actual_tr);
      end else begin
        `uvm_info("SCB", $sformatf("Actual: %s", actual_tr.convert2string()), UVM_MEDIUM)
      end
    end
  endtask
  
  //----------------------------------------------------------------------------
  // Compare with Expected Transaction
  //----------------------------------------------------------------------------
  function void compare_with_expected(i2c_transaction actual);
    i2c_transaction expected;
    bit matched = 1;
    
    // Get expected from queue
    expected = expected_queue.pop_front();
    total_compared++;
    
    // Compare address
    if (expected.addr !== actual.addr) begin
      matched = 0;
      `uvm_error("SCB", $sformatf("Address mismatch: exp=0x%02h, act=0x%02h",
                                  expected.addr, actual.addr))
    end
    
    // Compare direction (R/W)
    if (expected.direction !== actual.direction) begin
      matched = 0;
      `uvm_error("SCB", $sformatf("Direction mismatch: exp=%s, act=%s",
                                  expected.direction.name(), actual.direction.name()))
    end
    
    // Compare data
    if (expected.data.size() != actual.data.size()) begin
      matched = 0;
      `uvm_error("SCB", $sformatf("Data size mismatch: exp=%0d, act=%0d",
                                  expected.data.size(), actual.data.size()))
    end else begin
      foreach (expected.data[i]) begin
        if (expected.data[i] !== actual.data[i]) begin
          matched = 0;
          `uvm_error("SCB", $sformatf("Data[%0d] mismatch: exp=0x%02h, act=0x%02h",
                                      i, expected.data[i], actual.data[i]))
        end
      end
    end
    
    // Update statistics
    if (matched) begin
      total_matched++;
      `uvm_info("SCB", $sformatf("Transaction #%0d MATCHED", total_compared), UVM_MEDIUM)
    end else begin
      total_mismatched++;
      mismatch_event.trigger(actual);
    end
    
    // Trigger completion event
    comparison_done_event.trigger();
  endfunction
  
  //----------------------------------------------------------------------------
  // Add Expected Transaction (called from test/sequence)
  //----------------------------------------------------------------------------
  function void add_expected(i2c_transaction tr);
    i2c_transaction tr_copy;
    tr_copy = i2c_transaction::type_id::create("expected_tr");
    tr_copy.copy(tr);
    expected_queue.push_back(tr_copy);
    `uvm_info("SCB", $sformatf("Added expected: %s (queue size=%0d)", 
              tr.convert2string(), expected_queue.size()), UVM_HIGH)
  endfunction
  
  //----------------------------------------------------------------------------
  // Check Phase
  //----------------------------------------------------------------------------
  function void check_phase(uvm_phase phase);
    super.check_phase(phase);
    
    if (expected_queue.size() > 0)
      `uvm_error("SCB", $sformatf("%0d expected transactions unmatched", expected_queue.size()))
  endfunction
  
  //----------------------------------------------------------------------------
  // Report Phase - Statistics
  //----------------------------------------------------------------------------
  function void report_phase(uvm_phase phase);
    real match_rate;
    super.report_phase(phase);
    
    match_rate = (total_compared > 0) ? (100.0 * total_matched / total_compared) : 100.0;
    
    `uvm_info("SCB", "╔════════════════════════════════════╗", UVM_NONE)
    `uvm_info("SCB", "║    SCOREBOARD STATISTICS           ║", UVM_NONE)
    `uvm_info("SCB", "╠════════════════════════════════════╣", UVM_NONE)
    `uvm_info("SCB", $sformatf("║ Received:    %8d             ║", total_received), UVM_NONE)
    `uvm_info("SCB", $sformatf("║ Compared:    %8d             ║", total_compared), UVM_NONE)
    `uvm_info("SCB", $sformatf("║ Matched:     %8d             ║", total_matched), UVM_NONE)
    `uvm_info("SCB", $sformatf("║ Mismatched:  %8d             ║", total_mismatched), UVM_NONE)
    `uvm_info("SCB", $sformatf("║ Match Rate:  %7.1f%%            ║", match_rate), UVM_NONE)
    `uvm_info("SCB", "╚════════════════════════════════════╝", UVM_NONE)
  endfunction
  
  //----------------------------------------------------------------------------
  // Utility: Wait for N comparisons
  //----------------------------------------------------------------------------
  task wait_for_comparisons(int count = 1);
    repeat(count) begin
      comparison_done_event.wait_trigger();
      comparison_done_event.reset();
    end
  endtask

endclass

`endif // I2C_SCOREBOARD_SV
